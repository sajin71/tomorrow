package fpu_misc is

  type FPU_CTRL is (unko);
  type comp_t is (fEQ, fLT);
  type FPU_OPER is (O_FADD, O_FSUB, O_FMUL, O_FDIV, O_FSQRT, O_FABS, O_FNEG, O_FROUND, O_FFLOOR, O_FRECIP, O_FCVTS);

end fpu_misc;
